class rohit;

int r;
int b
endclass
