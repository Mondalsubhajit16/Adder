interface axi_if;
	logic resetn;
	logic ip1;
	logic ip2;
	logic out;
endinterface
